magic
tech sky130A
timestamp 1615382711
<< nwell >>
rect -107 -3 156 195
<< mvnmos >>
rect -21 -95 38 -43
<< mvpmos >>
rect -21 30 38 120
<< mvndiff >>
rect -72 -57 -21 -43
rect -72 -85 -60 -57
rect -36 -85 -21 -57
rect -72 -95 -21 -85
rect 38 -53 90 -43
rect 38 -79 50 -53
rect 67 -79 90 -53
rect 38 -95 90 -79
<< mvpdiff >>
rect -72 93 -21 120
rect -72 62 -59 93
rect -42 62 -21 93
rect -72 30 -21 62
rect 38 94 91 120
rect 38 63 50 94
rect 67 63 91 94
rect 38 30 91 63
<< mvndiffc >>
rect -60 -85 -36 -57
rect 50 -79 67 -53
<< mvpdiffc >>
rect -59 62 -42 93
rect 50 63 67 94
<< poly >>
rect -21 120 38 133
rect -21 -43 38 30
rect -21 -114 38 -95
<< locali >>
rect -64 188 -30 191
rect -92 182 144 188
rect -92 153 -68 182
rect -38 153 144 182
rect -92 149 144 153
rect -64 93 -30 149
rect -64 62 -59 93
rect -42 62 -30 93
rect -64 30 -30 62
rect 46 94 68 120
rect 46 63 50 94
rect 67 63 68 94
rect -64 -57 -30 -43
rect -64 -85 -60 -57
rect -36 -85 -30 -57
rect -64 -121 -30 -85
rect 46 -53 68 63
rect 46 -79 50 -53
rect 67 -79 68 -53
rect 46 -95 68 -79
rect -64 -124 90 -121
rect -64 -153 -61 -124
rect -31 -153 90 -124
rect -64 -155 90 -153
rect -64 -156 -30 -155
<< viali >>
rect -68 153 -38 182
rect -61 -153 -31 -124
<< metal1 >>
rect -97 182 147 191
rect -97 153 -68 182
rect -38 153 147 182
rect -97 144 147 153
rect -75 -124 94 -120
rect -75 -153 -61 -124
rect -31 -153 94 -124
rect -75 -156 94 -153
rect -48 -157 94 -156
<< end >>
