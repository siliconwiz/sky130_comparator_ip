magic
tech sky130A
timestamp 1614994375
<< nwell >>
rect -107 -3 156 195
<< nmos >>
rect -21 -95 38 -43
<< mvpmos >>
rect -21 30 38 120
<< ndiff >>
rect -72 -54 -21 -43
rect -72 -82 -58 -54
rect -41 -82 -21 -54
rect -72 -95 -21 -82
rect 38 -54 75 -43
rect 38 -82 49 -54
rect 66 -82 75 -54
rect 38 -95 75 -82
<< mvpdiff >>
rect -72 93 -21 120
rect -72 62 -59 93
rect -42 62 -21 93
rect -72 30 -21 62
rect 38 94 91 120
rect 38 63 50 94
rect 67 63 91 94
rect 38 30 91 63
<< ndiffc >>
rect -58 -82 -41 -54
rect 49 -82 66 -54
<< mvpdiffc >>
rect -59 62 -42 93
rect 50 63 67 94
<< poly >>
rect -21 120 38 133
rect -21 -43 38 30
rect -21 -114 38 -95
<< locali >>
rect -64 188 -30 191
rect -92 182 144 188
rect -92 153 -68 182
rect -38 153 144 182
rect -92 149 144 153
rect -64 93 -30 149
rect -64 62 -59 93
rect -42 62 -30 93
rect -64 30 -30 62
rect 46 94 68 120
rect 46 63 50 94
rect 67 63 68 94
rect -64 -54 -30 -42
rect -64 -82 -58 -54
rect -41 -82 -30 -54
rect -64 -121 -30 -82
rect 46 -54 68 63
rect 46 -82 49 -54
rect 66 -82 68 -54
rect 46 -95 68 -82
rect -64 -124 90 -121
rect -64 -153 -61 -124
rect -31 -153 90 -124
rect -64 -155 90 -153
rect -64 -156 -30 -155
<< viali >>
rect -68 153 -38 182
rect -61 -153 -31 -124
<< metal1 >>
rect -97 182 147 191
rect -97 153 -68 182
rect -38 153 147 182
rect -97 144 147 153
rect -75 -124 94 -120
rect -75 -153 -61 -124
rect -31 -153 94 -124
rect -75 -156 94 -153
rect -48 -157 94 -156
<< end >>
