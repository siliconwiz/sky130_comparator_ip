magic
tech sky130A
timestamp 1615603199
<< nwell >>
rect -210 100 782 800
<< mvnmos >>
rect -136 -150 -86 50
rect 33 -150 83 50
rect 173 -149 223 51z
rect 305 -150 355 50
rect 445 -150 495 50
rect 549 -150 599 50
rect 662 -150 712 50
rect 33 -410 83 -210
rect 173 -410 223 -210
rect 305 -410 355 -211
rect 445 -410 495 -210
<< mvpmos >>
rect -152 135 -52 235
rect -6 135 94 235
rect 305 135 355 735
rect 445 135 495 587
rect 549 135 599 587
rect 662 135 712 587
<< mvndiff >>
rect -179 -150 -136 50
rect -86 -150 33 50
rect 83 -150 118 50
rect 148 -149 173 51
rect 223 -149 249 51
rect 280 -150 305 50
rect 355 -150 383 50
rect 417 -150 445 50
rect 495 -150 549 50
rect 599 -150 662 50
rect 712 -150 747 50
rect -1 -410 33 -210
rect 83 -410 173 -210
rect 223 -410 249 -210
rect 417 -211 445 -210
rect 279 -410 305 -211
rect 355 -410 445 -211
rect 495 -410 530 -210
<< mvpdiff >>
rect -177 135 -152 235
rect -52 135 -6 235
rect 94 135 131 235
rect 278 135 305 735
rect 355 535 405 735
rect 355 135 445 535
rect 495 135 549 535
rect 599 135 662 535
rect 712 135 747 535
<< poly >>
rect 305 735 355 750
rect -152 235 -52 262
rect -6 235 94 262
rect -152 113 -52 135
rect -6 112 94 135
rect -136 50 -86 73
rect 33 50 83 73
rect 173 51 223 74
rect 305 50 355 135
rect 445 50 495 135
rect 549 50 599 135
rect 662 50 712 135
rect -136 -164 -86 -150
rect 33 -164 83 -150
rect 33 -210 83 -186
rect 173 -210 223 -149
rect 305 -164 355 -150
rect 445 -164 495 -150
rect 549 -164 599 -150
rect 662 -164 712 -150
rect 305 -211 355 -186
rect 445 -210 495 -186
rect 33 -441 83 -410
rect 173 -440 223 -410
rect 305 -441 355 -410
rect 445 -441 495 -410
<< end >>
