magic
tech sky130A
timestamp 1615801552
<< nwell >>
rect -243 102 799 810
rect -243 100 243 102
rect 445 100 799 102
<< mvnmos >>
rect -136 -114 -86 -14
rect 33 -114 83 -14
rect 257 -100 307 -50
rect 445 -214 495 -14
rect 549 -214 599 -14
rect 662 -214 712 -14
rect 131 -285 181 -235
rect -9 -403 91 -353
rect 131 -403 181 -353
rect 305 -568 355 -368
rect 445 -568 495 -368
<< mvpmos >>
rect -152 135 -52 235
rect -6 135 94 235
rect 257 135 307 735
rect 445 135 495 535
rect 549 135 599 535
rect 662 135 712 535
<< mvndiff >>
rect -208 -22 -136 -14
rect -208 -106 -191 -22
rect -162 -106 -136 -22
rect -208 -114 -136 -106
rect -86 -22 33 -14
rect -86 -106 -71 -22
rect 17 -106 33 -22
rect -86 -114 33 -106
rect 83 -22 153 -14
rect 83 -106 102 -22
rect 145 -106 153 -22
rect 405 -22 445 -14
rect 198 -58 257 -50
rect 198 -92 206 -58
rect 235 -92 257 -58
rect 198 -100 257 -92
rect 307 -58 349 -50
rect 307 -92 323 -58
rect 341 -92 349 -58
rect 307 -100 349 -92
rect 83 -114 153 -106
rect 405 -206 413 -22
rect 431 -206 445 -22
rect 405 -214 445 -206
rect 495 -214 549 -14
rect 599 -22 662 -14
rect 599 -206 616 -22
rect 644 -206 662 -22
rect 599 -214 662 -206
rect 712 -22 756 -14
rect 712 -206 727 -22
rect 748 -206 756 -22
rect 712 -214 756 -206
rect 97 -243 131 -235
rect 97 -277 102 -243
rect 119 -277 131 -243
rect 97 -285 131 -277
rect 181 -246 234 -235
rect 181 -275 202 -246
rect 228 -275 234 -246
rect 181 -285 234 -275
rect -57 -362 -9 -353
rect -57 -394 -48 -362
rect -26 -394 -9 -362
rect -57 -403 -9 -394
rect 91 -361 131 -353
rect 91 -395 102 -361
rect 119 -395 131 -361
rect 91 -403 131 -395
rect 181 -361 221 -353
rect 181 -395 194 -361
rect 213 -395 221 -361
rect 181 -403 221 -395
rect 258 -376 305 -368
rect 258 -557 269 -376
rect 295 -557 305 -376
rect 258 -568 305 -557
rect 355 -376 445 -368
rect 355 -560 372 -376
rect 430 -560 445 -376
rect 355 -568 445 -560
rect 495 -376 538 -368
rect 495 -560 510 -376
rect 530 -560 538 -376
rect 495 -568 538 -560
<< mvpdiff >>
rect 204 727 257 735
rect -206 228 -152 235
rect -206 143 -194 228
rect -176 143 -152 228
rect -206 135 -152 143
rect -52 227 -6 235
rect -52 144 -43 227
rect -15 144 -6 227
rect -52 135 -6 144
rect 94 227 153 235
rect 94 143 117 227
rect 145 143 153 227
rect 94 135 153 143
rect 204 143 212 727
rect 241 143 257 727
rect 204 135 257 143
rect 307 727 433 735
rect 307 143 322 727
rect 425 535 433 727
rect 425 143 445 535
rect 307 135 445 143
rect 495 527 549 535
rect 495 143 512 527
rect 532 143 549 527
rect 495 135 549 143
rect 599 527 662 535
rect 599 142 612 527
rect 648 142 662 527
rect 599 135 662 142
rect 712 527 756 535
rect 712 143 727 527
rect 748 143 756 527
rect 712 135 756 143
<< mvndiffc >>
rect -191 -106 -162 -22
rect -71 -106 17 -22
rect 102 -106 145 -22
rect 206 -92 235 -58
rect 323 -92 341 -58
rect 413 -206 431 -22
rect 616 -206 644 -22
rect 727 -206 748 -22
rect 102 -277 119 -243
rect 202 -275 228 -246
rect -48 -394 -26 -362
rect 102 -395 119 -361
rect 194 -395 213 -361
rect 269 -557 295 -376
rect 372 -560 430 -376
rect 510 -560 530 -376
<< mvpdiffc >>
rect -194 143 -176 228
rect -43 144 -15 227
rect 117 143 145 227
rect 212 143 241 727
rect 322 143 425 727
rect 512 143 532 527
rect 612 142 648 527
rect 727 143 748 527
<< poly >>
rect 257 735 307 750
rect -152 235 -52 262
rect -6 235 94 262
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 445 535 495 558
rect 549 535 599 566
rect 662 535 712 558
rect -152 110 -52 135
rect -152 93 -144 110
rect -59 93 -52 110
rect -152 85 -52 93
rect -6 110 94 135
rect -6 93 2 110
rect 87 93 94 110
rect -6 85 94 93
rect 257 110 307 135
rect 257 88 265 110
rect 299 88 307 110
rect 257 80 307 88
rect 445 110 495 135
rect 445 49 453 110
rect 487 49 495 110
rect 257 19 307 27
rect -136 -14 -86 -1
rect 33 -14 83 -1
rect 257 -12 266 19
rect 299 -12 307 19
rect 257 -50 307 -12
rect 445 -14 495 49
rect 549 -14 599 135
rect 662 106 712 135
rect 662 12 670 106
rect 704 12 712 106
rect 662 -14 712 12
rect 257 -113 307 -100
rect -136 -201 -86 -114
rect 33 -132 83 -114
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect -136 -239 -86 -231
rect 131 -235 181 -212
rect 445 -227 495 -214
rect 549 -227 599 -214
rect 662 -228 712 -214
rect 131 -310 181 -285
rect -9 -353 91 -329
rect 131 -330 139 -310
rect 173 -330 181 -310
rect 131 -353 181 -330
rect 445 -303 495 -295
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 305 -368 355 -344
rect 445 -368 495 -343
rect -9 -428 91 -403
rect -9 -457 -1 -428
rect 71 -457 91 -428
rect 131 -436 181 -403
rect -9 -465 91 -457
rect 305 -593 355 -568
rect 445 -583 495 -568
rect 305 -618 313 -593
rect 347 -618 355 -593
rect 305 -627 355 -618
<< polycont >>
rect 557 566 591 596
rect -144 93 -59 110
rect 2 93 87 110
rect 265 88 299 110
rect 453 49 487 110
rect 266 -12 299 19
rect 670 12 704 106
rect 41 -170 71 -140
rect -128 -231 -94 -201
rect 139 -330 173 -310
rect 453 -343 487 -303
rect -1 -457 71 -428
rect 313 -618 347 -593
<< locali >>
rect 250 798 799 810
rect 250 765 262 798
rect 293 765 799 798
rect 250 758 799 765
rect 204 727 249 735
rect -202 228 -167 235
rect -202 143 -194 228
rect -176 143 -167 228
rect -202 135 -167 143
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 109 227 153 235
rect 109 143 117 227
rect 145 143 153 227
rect 109 135 153 143
rect 204 143 212 727
rect 241 143 249 727
rect 204 135 249 143
rect 314 727 433 735
rect 314 143 322 727
rect 425 143 433 727
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 143
rect 504 527 540 535
rect 504 143 512 527
rect 532 143 540 527
rect 504 135 540 143
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 719 527 756 535
rect 719 143 727 527
rect 748 143 756 527
rect 719 135 756 143
rect -152 110 94 118
rect -152 93 -144 110
rect -59 93 2 110
rect 87 93 94 110
rect -152 85 94 93
rect 257 110 307 118
rect 257 88 265 110
rect 299 88 307 110
rect 257 80 307 88
rect 445 110 495 118
rect 445 49 453 110
rect 487 49 495 110
rect 445 41 495 49
rect 662 106 712 114
rect 257 19 307 27
rect 257 -12 266 19
rect 299 -12 307 19
rect 662 12 670 106
rect 704 12 712 106
rect 662 4 712 12
rect -203 -22 -148 -14
rect -203 -106 -191 -22
rect -162 -106 -148 -22
rect -203 -114 -148 -106
rect -79 -22 25 -14
rect -79 -106 -71 -22
rect 17 -106 25 -22
rect -79 -114 25 -106
rect 94 -22 153 -14
rect 257 -20 307 -12
rect 94 -106 102 -22
rect 145 -106 153 -22
rect 405 -22 439 -14
rect 198 -58 243 -50
rect 198 -92 206 -58
rect 235 -92 243 -58
rect 198 -100 243 -92
rect 315 -58 349 -50
rect 315 -92 323 -58
rect 341 -92 349 -58
rect 315 -100 349 -92
rect 94 -114 153 -106
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -201 -86 -193
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect 405 -206 413 -22
rect 431 -206 439 -22
rect 405 -214 439 -206
rect 608 -22 652 -14
rect 608 -206 616 -22
rect 644 -206 652 -22
rect 608 -214 652 -206
rect 719 -22 756 -14
rect 719 -206 727 -22
rect 748 -206 756 -22
rect 719 -214 756 -206
rect -136 -239 -86 -231
rect 97 -243 125 -235
rect 97 -277 102 -243
rect 119 -277 125 -243
rect 97 -285 125 -277
rect 185 -246 234 -235
rect 185 -275 202 -246
rect 228 -275 234 -246
rect 185 -285 234 -275
rect 185 -302 221 -285
rect 131 -310 221 -302
rect 131 -330 139 -310
rect 173 -330 221 -310
rect 131 -336 221 -330
rect 445 -303 495 -295
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect -57 -362 -17 -353
rect -57 -394 -48 -362
rect -26 -394 -17 -362
rect -57 -403 -17 -394
rect 97 -361 126 -353
rect 97 -395 102 -361
rect 119 -395 126 -361
rect -9 -428 79 -420
rect -9 -457 -1 -428
rect 71 -457 79 -428
rect -9 -465 79 -457
rect 97 -647 126 -395
rect 186 -361 221 -353
rect 186 -395 194 -361
rect 213 -395 221 -361
rect 186 -403 221 -395
rect 258 -376 305 -368
rect 258 -557 269 -376
rect 295 -557 305 -376
rect 258 -568 305 -557
rect 363 -376 438 -368
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
rect 503 -376 538 -368
rect 503 -560 510 -376
rect 530 -560 538 -376
rect 503 -568 538 -560
rect 305 -593 355 -585
rect 305 -618 313 -593
rect 347 -618 355 -593
rect 305 -627 355 -618
rect -232 -659 767 -647
rect -232 -697 -219 -659
rect -191 -697 -162 -659
rect -134 -697 -99 -659
rect -71 -697 767 -659
rect -232 -705 767 -697
<< viali >>
rect 262 765 293 798
rect -194 143 -176 228
rect -43 144 -15 227
rect 117 143 145 227
rect 212 143 241 727
rect 322 143 425 727
rect 557 566 591 596
rect 512 143 532 527
rect 612 142 648 527
rect 727 143 748 527
rect -144 93 -59 110
rect 2 93 87 110
rect 265 88 299 110
rect 453 49 487 110
rect 266 -12 299 19
rect 670 12 704 106
rect -191 -106 -162 -22
rect -71 -106 17 -22
rect 102 -106 145 -22
rect 206 -92 235 -58
rect 323 -92 341 -58
rect 41 -170 71 -140
rect -128 -231 -94 -201
rect 413 -206 431 -22
rect 616 -206 644 -22
rect 727 -206 748 -22
rect 102 -277 119 -243
rect 202 -275 228 -246
rect 453 -343 487 -303
rect -48 -394 -26 -362
rect 102 -395 119 -361
rect -1 -457 71 -428
rect 194 -395 213 -361
rect 269 -557 295 -376
rect 372 -560 430 -376
rect 510 -560 530 -376
rect 313 -618 347 -593
rect -219 -697 -191 -659
rect -162 -697 -134 -659
rect -99 -697 -71 -659
<< metal1 >>
rect 250 798 799 810
rect 250 765 262 798
rect 293 765 799 798
rect 250 758 799 765
rect 204 727 249 735
rect -203 228 -167 235
rect -203 143 -194 228
rect -176 143 -167 228
rect -203 118 -167 143
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 109 227 153 235
rect 109 143 117 227
rect 145 143 153 227
rect -203 110 94 118
rect -203 93 -144 110
rect -59 93 2 110
rect 87 93 94 110
rect -203 85 94 93
rect 109 117 153 143
rect 204 143 212 727
rect 241 143 249 727
rect 204 135 249 143
rect 314 727 433 735
rect 314 143 322 727
rect 425 143 433 727
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 143
rect 504 527 541 535
rect 504 143 512 527
rect 532 143 541 527
rect 504 135 541 143
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 719 527 756 535
rect 719 143 727 527
rect 748 143 756 527
rect 719 135 756 143
rect 109 110 388 117
rect 109 88 265 110
rect 299 88 388 110
rect -203 -22 -148 85
rect 109 80 388 88
rect 109 -14 153 80
rect -203 -106 -191 -22
rect -162 -106 -148 -22
rect -203 -114 -148 -106
rect -79 -22 25 -14
rect -79 -106 -71 -22
rect 17 -106 25 -22
rect -79 -114 25 -106
rect 94 -22 153 -14
rect 263 19 307 27
rect 263 -12 266 19
rect 299 -12 307 19
rect 263 -20 307 -12
rect 94 -106 102 -22
rect 145 -106 153 -22
rect 198 -58 243 -50
rect 198 -92 206 -58
rect 235 -92 243 -58
rect 198 -100 243 -92
rect 315 -58 349 -50
rect 315 -92 323 -58
rect 341 -92 349 -58
rect 94 -114 153 -106
rect -203 -528 -151 -114
rect -136 -201 -86 -193
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect -136 -239 -86 -231
rect -57 -362 -15 -114
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 33 -178 80 -170
rect 315 -182 349 -92
rect -57 -394 -48 -362
rect -26 -394 -15 -362
rect -57 -403 -15 -394
rect 97 -211 349 -182
rect 97 -243 126 -211
rect 97 -277 102 -243
rect 119 -277 126 -243
rect 97 -361 126 -277
rect 196 -246 234 -240
rect 196 -275 202 -246
rect 228 -275 234 -246
rect 196 -281 234 -275
rect 363 -263 388 80
rect 445 110 495 118
rect 445 49 453 110
rect 487 49 495 110
rect 445 41 495 49
rect 509 114 541 135
rect 509 106 712 114
rect 509 14 670 106
rect 405 12 670 14
rect 704 12 712 106
rect 405 4 712 12
rect 405 -14 541 4
rect 727 -14 756 135
rect 405 -22 439 -14
rect 405 -206 413 -22
rect 431 -206 439 -22
rect 405 -228 439 -206
rect 608 -22 652 -14
rect 608 -206 616 -22
rect 644 -206 652 -22
rect 405 -249 589 -228
rect 363 -279 538 -263
rect 445 -303 495 -295
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect 97 -395 102 -361
rect 119 -395 126 -361
rect 97 -403 126 -395
rect 186 -361 221 -353
rect 186 -395 194 -361
rect 220 -395 221 -361
rect 509 -368 538 -279
rect 186 -403 221 -395
rect 258 -376 305 -368
rect -9 -428 79 -420
rect -9 -457 -1 -428
rect 71 -457 79 -428
rect -9 -465 79 -457
rect 258 -528 269 -376
rect -203 -557 269 -528
rect 295 -557 305 -376
rect -203 -568 305 -557
rect 363 -376 438 -368
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
rect 503 -376 538 -368
rect 503 -560 510 -376
rect 530 -560 538 -376
rect 503 -568 538 -560
rect 561 -585 589 -249
rect 305 -593 591 -585
rect 305 -618 313 -593
rect 347 -618 591 -593
rect 305 -627 591 -618
rect 608 -647 652 -206
rect 719 -22 756 -14
rect 719 -206 727 -22
rect 748 -206 756 -22
rect 719 -214 756 -206
rect -232 -659 767 -647
rect -232 -697 -219 -659
rect -191 -697 -162 -659
rect -134 -697 -99 -659
rect -71 -697 767 -659
rect -232 -705 767 -697
<< via1 >>
rect 262 765 293 798
rect -43 144 -15 227
rect 322 143 425 727
rect 557 566 591 596
rect 612 142 648 527
rect 266 -12 299 19
rect -128 -231 -94 -201
rect 41 -170 71 -140
rect 202 -275 228 -246
rect 453 49 487 110
rect 453 -343 487 -303
rect 194 -395 213 -361
rect 213 -395 220 -361
rect -1 -457 71 -428
rect 372 -560 430 -376
<< metal2 >>
rect 250 798 799 810
rect 250 765 262 798
rect 293 765 799 798
rect 250 758 799 765
rect 314 727 433 735
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 314 143 322 727
rect 425 143 433 727
rect 549 603 846 648
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 143
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 204 72 243 135
rect 445 110 495 118
rect 445 72 453 110
rect 204 49 453 72
rect 487 49 495 110
rect 204 41 495 49
rect 204 -50 243 41
rect 257 19 307 27
rect 257 -12 266 19
rect 299 -12 307 19
rect 257 -20 307 -12
rect 198 -58 243 -50
rect 198 -92 206 -58
rect 235 -92 243 -58
rect 198 -100 243 -92
rect -275 -140 80 -132
rect -275 -170 41 -140
rect 71 -170 80 -140
rect -275 -178 80 -170
rect -361 -201 -86 -193
rect -361 -231 -128 -201
rect -94 -231 -86 -201
rect -361 -239 -86 -231
rect 196 -246 796 -235
rect 196 -275 202 -246
rect 228 -275 796 -246
rect 196 -281 796 -275
rect 196 -285 234 -281
rect 445 -303 495 -295
rect 221 -343 431 -319
rect 221 -353 250 -343
rect 186 -361 250 -353
rect 186 -395 194 -361
rect 220 -395 250 -361
rect 186 -403 250 -395
rect 363 -368 431 -343
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect 363 -376 438 -368
rect -9 -428 79 -420
rect -9 -457 -1 -428
rect 71 -457 79 -428
rect -9 -465 79 -457
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
<< via2 >>
rect -43 144 -15 227
rect 322 143 425 727
rect 612 142 648 527
rect 266 -12 299 19
rect 206 -92 235 -58
rect 453 -343 487 -303
rect -1 -457 71 -428
<< metal3 >>
rect -261 758 799 810
rect -261 -420 -226 758
rect -48 227 -10 758
rect 156 757 200 758
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 314 727 433 758
rect 314 143 322 727
rect 425 143 433 727
rect 314 135 433 143
rect 604 527 656 758
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 314 27 353 135
rect 257 19 353 27
rect 257 -12 266 19
rect 299 -12 353 19
rect 257 -20 353 -12
rect 198 -58 243 -50
rect 198 -92 206 -58
rect 235 -92 243 -58
rect 198 -125 243 -92
rect 198 -165 378 -125
rect 338 -295 378 -165
rect 338 -303 495 -295
rect 338 -338 453 -303
rect 445 -343 453 -338
rect 487 -343 495 -303
rect 445 -351 495 -343
rect -261 -428 79 -420
rect -261 -457 -1 -428
rect 71 -457 79 -428
rect -261 -465 79 -457
<< labels >>
rlabel metal1 159 -678 159 -678 1 GND
rlabel metal3 150 783 150 783 1 VDD
rlabel metal2 816 632 816 632 1 EN
rlabel metal2 759 -262 759 -262 1 Ihyst
rlabel metal2 -340 -224 -340 -224 1 INN
rlabel metal2 -271 -159 -271 -159 1 INP
<< end >>
